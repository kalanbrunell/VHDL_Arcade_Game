library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity thirtyTwoBlockROM is 
	port(
		clk : in std_logic;
		rowIn : in unsigned(9 downto 0);
		colIn : in unsigned(9 downto 0);
		rowOffset : in unsigned (9 downto 0);
		colOffset : in unsigned (9 downto 0);
		rgbOut : out std_logic_vector(5 downto 0)
	);
end;

architecture synth of thirtyTwoBlockROM is
	
	signal address : std_logic_vector(19 downto 0);
	signal offsetRow : unsigned(9 downto 0);
	signal offsetCol : unsigned(9 downto 0);
	signal scaleOffsetRow : unsigned(9 downto 0);
	signal scaleOffsetCol : unsigned(9 downto 0);
	signal rgb : std_logic_vector(5 downto 0);
	
	begin
		process(clk) begin
			if (rising_edge(clk)) then
				case address is
                    when "00000000000000000000" => rgb <= "100000";
                    when "00000000000000000001" => rgb <= "100000";
                    when "00000000000000000010" => rgb <= "100000";
                    when "00000000000000000011" => rgb <= "100000";
                    when "00000000000000000100" => rgb <= "100000";
                    when "00000000000000000101" => rgb <= "100000";
                    when "00000000000000000110" => rgb <= "100000";
                    when "00000000000000000111" => rgb <= "100000";
                    when "00000000000000001000" => rgb <= "100000";
                    when "00000000000000001001" => rgb <= "100000";
                    when "00000000000000001010" => rgb <= "100000";
                    when "00000000000000001011" => rgb <= "100000";
                    when "00000000000000001100" => rgb <= "100000";
                    when "00000000000000001101" => rgb <= "100000";
                    when "00000000000000001110" => rgb <= "100000";
                    when "00000000000000001111" => rgb <= "100000";
                    when "00000000010000000000" => rgb <= "100000";
                    when "00000000010000000001" => rgb <= "100000";
                    when "00000000010000000010" => rgb <= "100000";
                    when "00000000010000000011" => rgb <= "100000";
                    when "00000000010000000100" => rgb <= "100000";
                    when "00000000010000000101" => rgb <= "100000";
                    when "00000000010000000110" => rgb <= "100000";
                    when "00000000010000000111" => rgb <= "100000";
                    when "00000000010000001000" => rgb <= "100000";
                    when "00000000010000001001" => rgb <= "100000";
                    when "00000000010000001010" => rgb <= "100000";
                    when "00000000010000001011" => rgb <= "100000";
                    when "00000000010000001100" => rgb <= "100000";
                    when "00000000010000001101" => rgb <= "100000";
                    when "00000000010000001110" => rgb <= "100000";
                    when "00000000010000001111" => rgb <= "100000";
                    when "00000000100000000000" => rgb <= "100000";
                    when "00000000100000000001" => rgb <= "100000";
                    when "00000000100000000010" => rgb <= "100000";
                    when "00000000100000000011" => rgb <= "100000";
                    when "00000000100000000100" => rgb <= "100000";
                    when "00000000100000000101" => rgb <= "100000";
                    when "00000000100000000110" => rgb <= "100000";
                    when "00000000100000000111" => rgb <= "100000";
                    when "00000000100000001000" => rgb <= "100000";
                    when "00000000100000001001" => rgb <= "100000";
                    when "00000000100000001010" => rgb <= "100000";
                    when "00000000100000001011" => rgb <= "100000";
                    when "00000000100000001100" => rgb <= "100000";
                    when "00000000100000001101" => rgb <= "100000";
                    when "00000000100000001110" => rgb <= "100000";
                    when "00000000100000001111" => rgb <= "100000";
                    when "00000000110000000000" => rgb <= "100000";
                    when "00000000110000000001" => rgb <= "100000";
                    when "00000000110000000010" => rgb <= "100000";
                    when "00000000110000000011" => rgb <= "000000";
                    when "00000000110000000100" => rgb <= "000000";
                    when "00000000110000000101" => rgb <= "000000";
                    when "00000000110000000110" => rgb <= "000000";
                    when "00000000110000000111" => rgb <= "100000";
                    when "00000000110000001000" => rgb <= "100000";
                    when "00000000110000001001" => rgb <= "000000";
                    when "00000000110000001010" => rgb <= "000000";
                    when "00000000110000001011" => rgb <= "000000";
                    when "00000000110000001100" => rgb <= "000000";
                    when "00000000110000001101" => rgb <= "100000";
                    when "00000000110000001110" => rgb <= "100000";
                    when "00000000110000001111" => rgb <= "100000";
                    when "00000001000000000000" => rgb <= "100000";
                    when "00000001000000000001" => rgb <= "100000";
                    when "00000001000000000010" => rgb <= "100000";
                    when "00000001000000000011" => rgb <= "100000";
                    when "00000001000000000100" => rgb <= "100000";
                    when "00000001000000000101" => rgb <= "100000";
                    when "00000001000000000110" => rgb <= "000000";
                    when "00000001000000000111" => rgb <= "100000";
                    when "00000001000000001000" => rgb <= "100000";
                    when "00000001000000001001" => rgb <= "100000";
                    when "00000001000000001010" => rgb <= "100000";
                    when "00000001000000001011" => rgb <= "100000";
                    when "00000001000000001100" => rgb <= "000000";
                    when "00000001000000001101" => rgb <= "100000";
                    when "00000001000000001110" => rgb <= "100000";
                    when "00000001000000001111" => rgb <= "100000";
                    when "00000001010000000000" => rgb <= "100000";
                    when "00000001010000000001" => rgb <= "100000";
                    when "00000001010000000010" => rgb <= "100000";
                    when "00000001010000000011" => rgb <= "100000";
                    when "00000001010000000100" => rgb <= "100000";
                    when "00000001010000000101" => rgb <= "100000";
                    when "00000001010000000110" => rgb <= "000000";
                    when "00000001010000000111" => rgb <= "100000";
                    when "00000001010000001000" => rgb <= "100000";
                    when "00000001010000001001" => rgb <= "100000";
                    when "00000001010000001010" => rgb <= "100000";
                    when "00000001010000001011" => rgb <= "100000";
                    when "00000001010000001100" => rgb <= "000000";
                    when "00000001010000001101" => rgb <= "100000";
                    when "00000001010000001110" => rgb <= "100000";
                    when "00000001010000001111" => rgb <= "100000";
                    when "00000001100000000000" => rgb <= "100000";
                    when "00000001100000000001" => rgb <= "100000";
                    when "00000001100000000010" => rgb <= "100000";
                    when "00000001100000000011" => rgb <= "100000";
                    when "00000001100000000100" => rgb <= "100000";
                    when "00000001100000000101" => rgb <= "100000";
                    when "00000001100000000110" => rgb <= "000000";
                    when "00000001100000000111" => rgb <= "100000";
                    when "00000001100000001000" => rgb <= "100000";
                    when "00000001100000001001" => rgb <= "100000";
                    when "00000001100000001010" => rgb <= "100000";
                    when "00000001100000001011" => rgb <= "100000";
                    when "00000001100000001100" => rgb <= "000000";
                    when "00000001100000001101" => rgb <= "100000";
                    when "00000001100000001110" => rgb <= "100000";
                    when "00000001100000001111" => rgb <= "100000";
                    when "00000001110000000000" => rgb <= "100000";
                    when "00000001110000000001" => rgb <= "100000";
                    when "00000001110000000010" => rgb <= "100000";
                    when "00000001110000000011" => rgb <= "000000";
                    when "00000001110000000100" => rgb <= "000000";
                    when "00000001110000000101" => rgb <= "000000";
                    when "00000001110000000110" => rgb <= "000000";
                    when "00000001110000000111" => rgb <= "100000";
                    when "00000001110000001000" => rgb <= "100000";
                    when "00000001110000001001" => rgb <= "000000";
                    when "00000001110000001010" => rgb <= "000000";
                    when "00000001110000001011" => rgb <= "000000";
                    when "00000001110000001100" => rgb <= "000000";
                    when "00000001110000001101" => rgb <= "100000";
                    when "00000001110000001110" => rgb <= "100000";
                    when "00000001110000001111" => rgb <= "100000";
                    when "00000010000000000000" => rgb <= "100000";
                    when "00000010000000000001" => rgb <= "100000";
                    when "00000010000000000010" => rgb <= "100000";
                    when "00000010000000000011" => rgb <= "100000";
                    when "00000010000000000100" => rgb <= "100000";
                    when "00000010000000000101" => rgb <= "100000";
                    when "00000010000000000110" => rgb <= "000000";
                    when "00000010000000000111" => rgb <= "100000";
                    when "00000010000000001000" => rgb <= "100000";
                    when "00000010000000001001" => rgb <= "000000";
                    when "00000010000000001010" => rgb <= "100000";
                    when "00000010000000001011" => rgb <= "100000";
                    when "00000010000000001100" => rgb <= "100000";
                    when "00000010000000001101" => rgb <= "100000";
                    when "00000010000000001110" => rgb <= "100000";
                    when "00000010000000001111" => rgb <= "100000";
                    when "00000010010000000000" => rgb <= "100000";
                    when "00000010010000000001" => rgb <= "100000";
                    when "00000010010000000010" => rgb <= "100000";
                    when "00000010010000000011" => rgb <= "100000";
                    when "00000010010000000100" => rgb <= "100000";
                    when "00000010010000000101" => rgb <= "100000";
                    when "00000010010000000110" => rgb <= "000000";
                    when "00000010010000000111" => rgb <= "100000";
                    when "00000010010000001000" => rgb <= "100000";
                    when "00000010010000001001" => rgb <= "000000";
                    when "00000010010000001010" => rgb <= "100000";
                    when "00000010010000001011" => rgb <= "100000";
                    when "00000010010000001100" => rgb <= "100000";
                    when "00000010010000001101" => rgb <= "100000";
                    when "00000010010000001110" => rgb <= "100000";
                    when "00000010010000001111" => rgb <= "100000";
                    when "00000010100000000000" => rgb <= "100000";
                    when "00000010100000000001" => rgb <= "100000";
                    when "00000010100000000010" => rgb <= "100000";
                    when "00000010100000000011" => rgb <= "100000";
                    when "00000010100000000100" => rgb <= "100000";
                    when "00000010100000000101" => rgb <= "100000";
                    when "00000010100000000110" => rgb <= "000000";
                    when "00000010100000000111" => rgb <= "100000";
                    when "00000010100000001000" => rgb <= "100000";
                    when "00000010100000001001" => rgb <= "000000";
                    when "00000010100000001010" => rgb <= "100000";
                    when "00000010100000001011" => rgb <= "100000";
                    when "00000010100000001100" => rgb <= "100000";
                    when "00000010100000001101" => rgb <= "100000";
                    when "00000010100000001110" => rgb <= "100000";
                    when "00000010100000001111" => rgb <= "100000";
                    when "00000010110000000000" => rgb <= "100000";
                    when "00000010110000000001" => rgb <= "100000";
                    when "00000010110000000010" => rgb <= "100000";
                    when "00000010110000000011" => rgb <= "000000";
                    when "00000010110000000100" => rgb <= "000000";
                    when "00000010110000000101" => rgb <= "000000";
                    when "00000010110000000110" => rgb <= "000000";
                    when "00000010110000000111" => rgb <= "100000";
                    when "00000010110000001000" => rgb <= "100000";
                    when "00000010110000001001" => rgb <= "000000";
                    when "00000010110000001010" => rgb <= "000000";
                    when "00000010110000001011" => rgb <= "000000";
                    when "00000010110000001100" => rgb <= "000000";
                    when "00000010110000001101" => rgb <= "100000";
                    when "00000010110000001110" => rgb <= "100000";
                    when "00000010110000001111" => rgb <= "100000";
                    when "00000011000000000000" => rgb <= "100000";
                    when "00000011000000000001" => rgb <= "100000";
                    when "00000011000000000010" => rgb <= "100000";
                    when "00000011000000000011" => rgb <= "100000";
                    when "00000011000000000100" => rgb <= "100000";
                    when "00000011000000000101" => rgb <= "100000";
                    when "00000011000000000110" => rgb <= "100000";
                    when "00000011000000000111" => rgb <= "100000";
                    when "00000011000000001000" => rgb <= "100000";
                    when "00000011000000001001" => rgb <= "100000";
                    when "00000011000000001010" => rgb <= "100000";
                    when "00000011000000001011" => rgb <= "100000";
                    when "00000011000000001100" => rgb <= "100000";
                    when "00000011000000001101" => rgb <= "100000";
                    when "00000011000000001110" => rgb <= "100000";
                    when "00000011000000001111" => rgb <= "100000";
                    when "00000011010000000000" => rgb <= "100000";
                    when "00000011010000000001" => rgb <= "100000";
                    when "00000011010000000010" => rgb <= "100000";
                    when "00000011010000000011" => rgb <= "100000";
                    when "00000011010000000100" => rgb <= "100000";
                    when "00000011010000000101" => rgb <= "100000";
                    when "00000011010000000110" => rgb <= "100000";
                    when "00000011010000000111" => rgb <= "100000";
                    when "00000011010000001000" => rgb <= "100000";
                    when "00000011010000001001" => rgb <= "100000";
                    when "00000011010000001010" => rgb <= "100000";
                    when "00000011010000001011" => rgb <= "100000";
                    when "00000011010000001100" => rgb <= "100000";
                    when "00000011010000001101" => rgb <= "100000";
                    when "00000011010000001110" => rgb <= "100000";
                    when "00000011010000001111" => rgb <= "100000";
                    when "00000011100000000000" => rgb <= "100000";
                    when "00000011100000000001" => rgb <= "100000";
                    when "00000011100000000010" => rgb <= "100000";
                    when "00000011100000000011" => rgb <= "100000";
                    when "00000011100000000100" => rgb <= "100000";
                    when "00000011100000000101" => rgb <= "100000";
                    when "00000011100000000110" => rgb <= "100000";
                    when "00000011100000000111" => rgb <= "100000";
                    when "00000011100000001000" => rgb <= "100000";
                    when "00000011100000001001" => rgb <= "100000";
                    when "00000011100000001010" => rgb <= "100000";
                    when "00000011100000001011" => rgb <= "100000";
                    when "00000011100000001100" => rgb <= "100000";
                    when "00000011100000001101" => rgb <= "100000";
                    when "00000011100000001110" => rgb <= "100000";
                    when "00000011100000001111" => rgb <= "100000";
                    when "00000011110000000000" => rgb <= "100000";
                    when "00000011110000000001" => rgb <= "100000";
                    when "00000011110000000010" => rgb <= "100000";
                    when "00000011110000000011" => rgb <= "100000";
                    when "00000011110000000100" => rgb <= "100000";
                    when "00000011110000000101" => rgb <= "100000";
                    when "00000011110000000110" => rgb <= "100000";
                    when "00000011110000000111" => rgb <= "100000";
                    when "00000011110000001000" => rgb <= "100000";
                    when "00000011110000001001" => rgb <= "100000";
                    when "00000011110000001010" => rgb <= "100000";
                    when "00000011110000001011" => rgb <= "100000";
                    when "00000011110000001100" => rgb <= "100000";
                    when "00000011110000001101" => rgb <= "100000";
                    when "00000011110000001110" => rgb <= "100000";
                    when "00000011110000001111" => rgb <= "100000";
                    when others => rgb <= "000000";
					end case;
			end if;
	end process;

	offsetRow <= rowIn - rowOffset;
	offsetCol <= colIn - colOffset;
	scaleOffsetRow <= offsetRow / 4;
	scaleOffsetCol <= offsetCol / 4;
	address <= std_logic_vector(scaleOffsetRow) & std_logic_vector(scaleOffsetCol);
	rgbOut <= rgb;
end;